module KeyExpansion
(
  key,
  expandedKey
);

  localparam NB = 4;
  localparam NK = 8; //can be 4 for AES 128, 6 for AES 192 and 8 for AES 256 :number of words in key
  //TODO: represent NR as a function of NK
  localparam NR = 14; //can be 10 for AES 128, 12 for AES 256, and 14 for AES 512 (NR = NK+6)

  //AES takes 128bit or 256bit key and generates NR+1 128-bit subkeys out of it
  //So subkeys for the rounds are ALWAYS 128bit
  input     [(NK*32)-1:0]          key;
  output    [((NB*32)*(NR+1))-1:0] expandedKey;
  // expanded key = of 4*Nb*(Nr+1) bytes

  wire      [31:0]           w[NK*(NR+1)-1:0]; //number of words, each being 32bit (4 bytes)
  wire      [31:0]           t[NR-1:0];
  wire      [31:0]           tt[4*(NR+1)-1:0];
  wire      [7:0]            RCon[13:0];
  wire      [31:0]           rotWord[NR-1:0];
  wire      [31:0]           Q[NR-1:0];
  wire      [95:0]           unused[NR-1:0];
  wire      [95:0]           unused2[4*(NR+1)-1:0];

  /*unsigned char rcon[256] = {
    0x8d, 0x01, 0x02, 0x04, 0x08, 0x10, 0x20, 0x40, 0x80, 0x1b, 0x36, 0x6c, 0xd8, 0xab, 0x4d, 0x9a, 
    0x2f, 0x5e, 0xbc, 0x63, 0xc6, 0x97, 0x35, 0x6a, 0xd4, 0xb3, 0x7d, 0xfa, 0xef, 0xc5, 0x91, 0x39, 
    0x72, 0xe4, 0xd3, 0xbd, 0x61, 0xc2, 0x9f, 0x25, 0x4a, 0x94, 0x33, 0x66, 0xcc, 0x83, 0x1d, 0x3a, 
    0x74, 0xe8, 0xcb, 0x8d, 0x01, 0x02, 0x04, 0x08, 0x10, 0x20, 0x40, 0x80, 0x1b, 0x36, 0x6c, 0xd8, 
    0xab, 0x4d, 0x9a, 0x2f, 0x5e, 0xbc, 0x63, 0xc6, 0x97, 0x35, 0x6a, 0xd4, 0xb3, 0x7d, 0xfa, 0xef, 
    0xc5, 0x91, 0x39, 0x72, 0xe4, 0xd3, 0xbd, 0x61, 0xc2, 0x9f, 0x25, 0x4a, 0x94, 0x33, 0x66, 0xcc, 
    0x83, 0x1d, 0x3a, 0x74, 0xe8, 0xcb, 0x8d, 0x01, 0x02, 0x04, 0x08, 0x10, 0x20, 0x40, 0x80, 0x1b, 
    0x36, 0x6c, 0xd8, 0xab, 0x4d, 0x9a, 0x2f, 0x5e, 0xbc, 0x63, 0xc6, 0x97, 0x35, 0x6a, 0xd4, 0xb3, 
    0x7d, 0xfa, 0xef, 0xc5, 0x91, 0x39, 0x72, 0xe4, 0xd3, 0xbd, 0x61, 0xc2, 0x9f, 0x25, 0x4a, 0x94, 
    0x33, 0x66, 0xcc, 0x83, 0x1d, 0x3a, 0x74, 0xe8, 0xcb, 0x8d, 0x01, 0x02, 0x04, 0x08, 0x10, 0x20, 
    0x40, 0x80, 0x1b, 0x36, 0x6c, 0xd8, 0xab, 0x4d, 0x9a, 0x2f, 0x5e, 0xbc, 0x63, 0xc6, 0x97, 0x35, 
    0x6a, 0xd4, 0xb3, 0x7d, 0xfa, 0xef, 0xc5, 0x91, 0x39, 0x72, 0xe4, 0xd3, 0xbd, 0x61, 0xc2, 0x9f, 
    0x25, 0x4a, 0x94, 0x33, 0x66, 0xcc, 0x83, 0x1d, 0x3a, 0x74, 0xe8, 0xcb, 0x8d, 0x01, 0x02, 0x04, 
    0x08, 0x10, 0x20, 0x40, 0x80, 0x1b, 0x36, 0x6c, 0xd8, 0xab, 0x4d, 0x9a, 0x2f, 0x5e, 0xbc, 0x63, 
    0xc6, 0x97, 0x35, 0x6a, 0xd4, 0xb3, 0x7d, 0xfa, 0xef, 0xc5, 0x91, 0x39, 0x72, 0xe4, 0xd3, 0xbd, 
    0x61, 0xc2, 0x9f, 0x25, 0x4a, 0x94, 0x33, 0x66, 0xcc, 0x83, 0x1d, 0x3a, 0x74, 0xe8, 0xcb, 0x8d
}*/
	
  // only need some of Rcon values, for AES 128 up to Rcon[10] of the origianl Rcon matrix
  // for AES 256 up to Rcon[14] of original Rcon matrix
  // each round requires Rcon value
  // rcon[0] is not used in AES algorithm

  assign RCon[0] = 8'h01;
  assign RCon[1] = 8'h02;
  assign RCon[2] = 8'h04;
  assign RCon[3] = 8'h08;
  assign RCon[4] = 8'h10;
  assign RCon[5] = 8'h20;
  assign RCon[6] = 8'h40;
  assign RCon[7] = 8'h80;
  assign RCon[8] = 8'h1b;
  assign RCon[9] = 8'h36;
  assign RCon[10] = 8'h6c;
  assign RCon[11] = 8'hd8;
  assign RCon[12] = 8'hab;
  assign RCon[13] = 8'h4d;
  
  genvar i;

  generate 
  for(i=0;i<NB*(NR+1);i=i+1) //number of words generated, for AES 256 = 60 words, each word is 4 bytes = 32 bits
  begin:EXPANDKEY
    assign expandedKey[32*(i+1)-1:32*i] = w[i]; //assign each word (32 bit) to the expanded key
  end
  endgenerate


  generate 
  for(i=0;i<NB*(NR+1);i=i+1) begin:NR_W
    if(i<NK) begin:INITIAL
      assign w[i] = key[32*(i+1)-1:32*i];
    end else begin:NEXT
      if(i%NK==0) begin:FIRST
        assign w[i] = w[i-NK] ^ t[i/NK-1];
      end else begin: NEXT
	if (NK > 6 && (i%NK) == 4)  begin:NEXT
	  assign w[i] = w[i-NK] ^ tt[i];
        end else begin
            assign w[i] = w[i-1] ^ w[i-NK];
 	end
      end
    end
  end
  endgenerate


  generate 
  for(i=0;i<NR;i=i+1) begin:COREKEY
    assign rotWord[i] = {w[NK+NK*i-1][7:0], w[NK+NK*i-1][31:8]}; //only for words which are multiples of NK
    SubBytes b(.x({rotWord[i], 96'b0}), .z({Q[i], unused[i]}));
    assign t[i] = {Q[i][31:8], RCon[i] ^ Q[i][7:0]};
  end
  endgenerate

 generate
 for (i = 0; i < NB*(NR+1); i=i+1) begin: SBOX_ONLY
	if (NK > 6 && (i%NK) == 4)  begin
	   SubBytes c(.x({w[i-1], 96'b0}), .z({tt[i], unused2[i]}));
	end
	
 end
 endgenerate



endmodule


